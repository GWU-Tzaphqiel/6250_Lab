`timescale 1ns/10ps
`define DELAY 5
