module tb_fulladd;

reg [1:0] a,b;
reg cin;
wire [1:0]s;
wire cout;
integer i;

fulladder_2b U0(
.a(a),
.b(b),
.cin(cin),
.cout(cout),
.s(s));

initial begin
	a <= 0;
	b <= 0;
	cin <= 0;
	
	for (i = 0; i < 25; i = i + 1) begin
		#10 a <= $random;
			b <= $random;
				cin <= $random;
	end
	$stop;
end
endmodule