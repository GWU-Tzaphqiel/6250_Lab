/home/ead/G34397914/cadence/innovus/osu05_stdcells.lef